/*Automatically generated by parse-opcodes */
`include "Opcodes.defines"
import RVTypes::*;

//typedef enum {
//    Gpr,
//    Fpu,
//    None
//} RegType deriving (Bits, Eq, FShow);
//
//typedef enum {
//    S,
//    SB,
//    U,
//    UJ,
//    I,
//    Z,
//    None
//} ImmType deriving (Bits, Eq, FShow);

typedef struct {
    Maybe#(RegType) rs1;
    Maybe#(RegType) rs2;
    Maybe#(RegType) rs3;
    Maybe#(RegType) dst;
    ImmType imm;
} InstType deriving (Bits, Eq, FShow);

function InstType toInstType(Instruction inst);
    Maybe#(RegType) i = tagged Valid Gpr;
    Maybe#(RegType) f = tagged Valid Fpu;
    Maybe#(RegType) _ = tagged Invalid;
    InstType ret = (case (inst) matches
            `BEQ:        InstType{rs1: i, rs2: i, rs3: _, dst: _, imm:   SB};
            `BNE:        InstType{rs1: i, rs2: i, rs3: _, dst: _, imm:   SB};
            `BLT:        InstType{rs1: i, rs2: i, rs3: _, dst: _, imm:   SB};
            `BGE:        InstType{rs1: i, rs2: i, rs3: _, dst: _, imm:   SB};
            `BLTU:       InstType{rs1: i, rs2: i, rs3: _, dst: _, imm:   SB};
            `BGEU:       InstType{rs1: i, rs2: i, rs3: _, dst: _, imm:   SB};
            `JALR:       InstType{rs1: i, rs2: _, rs3: _, dst: i, imm:    I};
            `JAL:        InstType{rs1: _, rs2: _, rs3: _, dst: i, imm:   UJ};
            `LUI:        InstType{rs1: _, rs2: _, rs3: _, dst: i, imm:    U};
            `AUIPC:      InstType{rs1: _, rs2: _, rs3: _, dst: i, imm:    U};
            `ADDI:       InstType{rs1: i, rs2: _, rs3: _, dst: i, imm:    I};
            `SLLI:       InstType{rs1: i, rs2: _, rs3: _, dst: i, imm:    I};
            `SLTI:       InstType{rs1: i, rs2: _, rs3: _, dst: i, imm:    I};
            `SLTIU:      InstType{rs1: i, rs2: _, rs3: _, dst: i, imm:    I};
            `XORI:       InstType{rs1: i, rs2: _, rs3: _, dst: i, imm:    I};
            `SRLI:       InstType{rs1: i, rs2: _, rs3: _, dst: i, imm:    I};
            `SRAI:       InstType{rs1: i, rs2: _, rs3: _, dst: i, imm:    I};
            `ORI:        InstType{rs1: i, rs2: _, rs3: _, dst: i, imm:    I};
            `ANDI:       InstType{rs1: i, rs2: _, rs3: _, dst: i, imm:    I};
            `ADD:        InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `SUB:        InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `SLL:        InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `SLT:        InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `SLTU:       InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `XOR:        InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `SRL:        InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `SRA:        InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `OR:         InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `AND:        InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `ADDIW:      InstType{rs1: i, rs2: _, rs3: _, dst: i, imm:    I};
            `SLLIW:      InstType{rs1: i, rs2: _, rs3: _, dst: i, imm:    I};
            `SRLIW:      InstType{rs1: i, rs2: _, rs3: _, dst: i, imm:    I};
            `SRAIW:      InstType{rs1: i, rs2: _, rs3: _, dst: i, imm:    I};
            `ADDW:       InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `SUBW:       InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `SLLW:       InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `SRLW:       InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `SRAW:       InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `LB:         InstType{rs1: i, rs2: _, rs3: _, dst: i, imm:    I};
            `LH:         InstType{rs1: i, rs2: _, rs3: _, dst: i, imm:    I};
            `LW:         InstType{rs1: i, rs2: _, rs3: _, dst: i, imm:    I};
            `LD:         InstType{rs1: i, rs2: _, rs3: _, dst: i, imm:    I};
            `LBU:        InstType{rs1: i, rs2: _, rs3: _, dst: i, imm:    I};
            `LHU:        InstType{rs1: i, rs2: _, rs3: _, dst: i, imm:    I};
            `LWU:        InstType{rs1: i, rs2: _, rs3: _, dst: i, imm:    I};
            `SB:         InstType{rs1: i, rs2: i, rs3: _, dst: _, imm:    S};
            `SH:         InstType{rs1: i, rs2: i, rs3: _, dst: _, imm:    S};
            `SW:         InstType{rs1: i, rs2: i, rs3: _, dst: _, imm:    S};
            `SD:         InstType{rs1: i, rs2: i, rs3: _, dst: _, imm:    S};
            `FENCE:      InstType{rs1: _, rs2: _, rs3: _, dst: _, imm: None};
            `FENCE_I:    InstType{rs1: _, rs2: _, rs3: _, dst: _, imm: None};
            `MUL:        InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `MULH:       InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `MULHSU:     InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `MULHU:      InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `DIV:        InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `DIVU:       InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `REM:        InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `REMU:       InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `MULW:       InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `DIVW:       InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `DIVUW:      InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `REMW:       InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `REMUW:      InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `AMOADD_W:   InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `AMOXOR_W:   InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `AMOOR_W:    InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `AMOAND_W:   InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `AMOMIN_W:   InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `AMOMAX_W:   InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `AMOMINU_W:  InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `AMOMAXU_W:  InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `AMOSWAP_W:  InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `LR_W:       InstType{rs1: i, rs2: _, rs3: _, dst: i, imm: None};
            `SC_W:       InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `AMOADD_D:   InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `AMOXOR_D:   InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `AMOOR_D:    InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `AMOAND_D:   InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `AMOMIN_D:   InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `AMOMAX_D:   InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `AMOMINU_D:  InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `AMOMAXU_D:  InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `AMOSWAP_D:  InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `LR_D:       InstType{rs1: i, rs2: _, rs3: _, dst: i, imm: None};
            `SC_D:       InstType{rs1: i, rs2: i, rs3: _, dst: i, imm: None};
            `SCALL:      InstType{rs1: _, rs2: _, rs3: _, dst: _, imm: None};
            `SBREAK:     InstType{rs1: _, rs2: _, rs3: _, dst: _, imm: None};
            `SRET:       InstType{rs1: _, rs2: _, rs3: _, dst: _, imm: None};
            `SFENCE_VM:  InstType{rs1: i, rs2: _, rs3: _, dst: _, imm: None};
            `WFI:        InstType{rs1: _, rs2: _, rs3: _, dst: _, imm: None};
            `MRTH:       InstType{rs1: _, rs2: _, rs3: _, dst: _, imm: None};
            `MRTS:       InstType{rs1: _, rs2: _, rs3: _, dst: _, imm: None};
            `HRTS:       InstType{rs1: _, rs2: _, rs3: _, dst: _, imm: None};
            `CSRRW:      InstType{rs1: i, rs2: _, rs3: _, dst: i, imm: None};
            `CSRRS:      InstType{rs1: i, rs2: _, rs3: _, dst: i, imm: None};
            `CSRRC:      InstType{rs1: i, rs2: _, rs3: _, dst: i, imm: None};
            `CSRRWI:     InstType{rs1: _, rs2: _, rs3: _, dst: i, imm:    Z};
            `CSRRSI:     InstType{rs1: _, rs2: _, rs3: _, dst: i, imm:    Z};
            `CSRRCI:     InstType{rs1: _, rs2: _, rs3: _, dst: i, imm:    Z};
            `FADD_S:     InstType{rs1: f, rs2: f, rs3: _, dst: f, imm: None};
            `FSUB_S:     InstType{rs1: f, rs2: f, rs3: _, dst: f, imm: None};
            `FMUL_S:     InstType{rs1: f, rs2: f, rs3: _, dst: f, imm: None};
            `FDIV_S:     InstType{rs1: f, rs2: f, rs3: _, dst: f, imm: None};
            `FSGNJ_S:    InstType{rs1: f, rs2: f, rs3: _, dst: f, imm: None};
            `FSGNJN_S:   InstType{rs1: f, rs2: f, rs3: _, dst: f, imm: None};
            `FSGNJX_S:   InstType{rs1: f, rs2: f, rs3: _, dst: f, imm: None};
            `FMIN_S:     InstType{rs1: f, rs2: f, rs3: _, dst: f, imm: None};
            `FMAX_S:     InstType{rs1: f, rs2: f, rs3: _, dst: f, imm: None};
            `FSQRT_S:    InstType{rs1: f, rs2: _, rs3: _, dst: f, imm: None};
            `FADD_D:     InstType{rs1: f, rs2: f, rs3: _, dst: f, imm: None};
            `FSUB_D:     InstType{rs1: f, rs2: f, rs3: _, dst: f, imm: None};
            `FMUL_D:     InstType{rs1: f, rs2: f, rs3: _, dst: f, imm: None};
            `FDIV_D:     InstType{rs1: f, rs2: f, rs3: _, dst: f, imm: None};
            `FSGNJ_D:    InstType{rs1: f, rs2: f, rs3: _, dst: f, imm: None};
            `FSGNJN_D:   InstType{rs1: f, rs2: f, rs3: _, dst: f, imm: None};
            `FSGNJX_D:   InstType{rs1: f, rs2: f, rs3: _, dst: f, imm: None};
            `FMIN_D:     InstType{rs1: f, rs2: f, rs3: _, dst: f, imm: None};
            `FMAX_D:     InstType{rs1: f, rs2: f, rs3: _, dst: f, imm: None};
            `FCVT_S_D:   InstType{rs1: f, rs2: _, rs3: _, dst: f, imm: None};
            `FCVT_D_S:   InstType{rs1: f, rs2: _, rs3: _, dst: f, imm: None};
            `FSQRT_D:    InstType{rs1: f, rs2: _, rs3: _, dst: f, imm: None};
            `FLE_S:      InstType{rs1: f, rs2: f, rs3: _, dst: i, imm: None};
            `FLT_S:      InstType{rs1: f, rs2: f, rs3: _, dst: i, imm: None};
            `FEQ_S:      InstType{rs1: f, rs2: f, rs3: _, dst: i, imm: None};
            `FLE_D:      InstType{rs1: f, rs2: f, rs3: _, dst: i, imm: None};
            `FLT_D:      InstType{rs1: f, rs2: f, rs3: _, dst: i, imm: None};
            `FEQ_D:      InstType{rs1: f, rs2: f, rs3: _, dst: i, imm: None};
            `FCVT_W_S:   InstType{rs1: f, rs2: _, rs3: _, dst: i, imm: None};
            `FCVT_WU_S:  InstType{rs1: f, rs2: _, rs3: _, dst: i, imm: None};
            `FCVT_L_S:   InstType{rs1: f, rs2: _, rs3: _, dst: i, imm: None};
            `FCVT_LU_S:  InstType{rs1: f, rs2: _, rs3: _, dst: i, imm: None};
            `FMV_X_S:    InstType{rs1: f, rs2: _, rs3: _, dst: i, imm: None};
            `FCLASS_S:   InstType{rs1: f, rs2: _, rs3: _, dst: i, imm: None};
            `FCVT_W_D:   InstType{rs1: f, rs2: _, rs3: _, dst: i, imm: None};
            `FCVT_WU_D:  InstType{rs1: f, rs2: _, rs3: _, dst: i, imm: None};
            `FCVT_L_D:   InstType{rs1: f, rs2: _, rs3: _, dst: i, imm: None};
            `FCVT_LU_D:  InstType{rs1: f, rs2: _, rs3: _, dst: i, imm: None};
            `FMV_X_D:    InstType{rs1: f, rs2: _, rs3: _, dst: i, imm: None};
            `FCLASS_D:   InstType{rs1: f, rs2: _, rs3: _, dst: i, imm: None};
            `FCVT_S_W:   InstType{rs1: i, rs2: _, rs3: _, dst: f, imm: None};
            `FCVT_S_WU:  InstType{rs1: i, rs2: _, rs3: _, dst: f, imm: None};
            `FCVT_S_L:   InstType{rs1: i, rs2: _, rs3: _, dst: f, imm: None};
            `FCVT_S_LU:  InstType{rs1: i, rs2: _, rs3: _, dst: f, imm: None};
            `FMV_S_X:    InstType{rs1: i, rs2: _, rs3: _, dst: f, imm: None};
            `FCVT_D_W:   InstType{rs1: i, rs2: _, rs3: _, dst: f, imm: None};
            `FCVT_D_WU:  InstType{rs1: i, rs2: _, rs3: _, dst: f, imm: None};
            `FCVT_D_L:   InstType{rs1: i, rs2: _, rs3: _, dst: f, imm: None};
            `FCVT_D_LU:  InstType{rs1: i, rs2: _, rs3: _, dst: f, imm: None};
            `FMV_D_X:    InstType{rs1: i, rs2: _, rs3: _, dst: f, imm: None};
            `FLW:        InstType{rs1: i, rs2: _, rs3: _, dst: f, imm:    I};
            `FLD:        InstType{rs1: i, rs2: _, rs3: _, dst: f, imm:    I};
            `FSW:        InstType{rs1: i, rs2: f, rs3: _, dst: _, imm:    S};
            `FSD:        InstType{rs1: i, rs2: f, rs3: _, dst: _, imm:    S};
            `FMADD_S:    InstType{rs1: f, rs2: f, rs3: f, dst: f, imm: None};
            `FMSUB_S:    InstType{rs1: f, rs2: f, rs3: f, dst: f, imm: None};
            `FNMSUB_S:   InstType{rs1: f, rs2: f, rs3: f, dst: f, imm: None};
            `FNMADD_S:   InstType{rs1: f, rs2: f, rs3: f, dst: f, imm: None};
            `FMADD_D:    InstType{rs1: f, rs2: f, rs3: f, dst: f, imm: None};
            `FMSUB_D:    InstType{rs1: f, rs2: f, rs3: f, dst: f, imm: None};
            `FNMSUB_D:   InstType{rs1: f, rs2: f, rs3: f, dst: f, imm: None};
            `FNMADD_D:   InstType{rs1: f, rs2: f, rs3: f, dst: f, imm: None};
            default:     ?;
        endcase);
    if ((ret.dst == tagged Valid Gpr) && (getInstFields(inst).rd == 0)) begin
        ret.dst = tagged Invalid;
    end
    return ret;
endfunction

//typedef enum {
//    CSRfflags       = 12'h001,
//    CSRfrm          = 12'h002,
//    CSRfcsr         = 12'h003,
//    CSRcycle        = 12'hc00,
//    CSRtime         = 12'hc01,
//    CSRinstret      = 12'hc02,
//    CSRstats        = 12'h0c0,
//    CSRuarch0       = 12'hcc0,
//    CSRuarch1       = 12'hcc1,
//    CSRuarch2       = 12'hcc2,
//    CSRuarch3       = 12'hcc3,
//    CSRuarch4       = 12'hcc4,
//    CSRuarch5       = 12'hcc5,
//    CSRuarch6       = 12'hcc6,
//    CSRuarch7       = 12'hcc7,
//    CSRuarch8       = 12'hcc8,
//    CSRuarch9       = 12'hcc9,
//    CSRuarch10      = 12'hcca,
//    CSRuarch11      = 12'hccb,
//    CSRuarch12      = 12'hccc,
//    CSRuarch13      = 12'hccd,
//    CSRuarch14      = 12'hcce,
//    CSRuarch15      = 12'hccf,
//    CSRsstatus      = 12'h100,
//    CSRstvec        = 12'h101,
//    CSRsie          = 12'h104,
//    CSRsscratch     = 12'h140,
//    CSRsepc         = 12'h141,
//    CSRsip          = 12'h144,
//    CSRsptbr        = 12'h180,
//    CSRsasid        = 12'h181,
//    CSRcyclew       = 12'h900,
//    CSRtimew        = 12'h901,
//    CSRinstretw     = 12'h902,
//    CSRstime        = 12'hd01,
//    CSRscause       = 12'hd42,
//    CSRsbadaddr     = 12'hd43,
//    CSRstimew       = 12'ha01,
//    CSRmstatus      = 12'h300,
//    CSRmtvec        = 12'h301,
//    CSRmtdeleg      = 12'h302,
//    CSRmie          = 12'h304,
//    CSRmtimecmp     = 12'h321,
//    CSRmscratch     = 12'h340,
//    CSRmepc         = 12'h341,
//    CSRmcause       = 12'h342,
//    CSRmbadaddr     = 12'h343,
//    CSRmip          = 12'h344,
//    CSRmtime        = 12'h701,
//    CSRmcpuid       = 12'hf00,
//    CSRmimpid       = 12'hf01,
//    CSRmhartid      = 12'hf10,
//    CSRmtohost      = 12'h780,
//    CSRmfromhost    = 12'h781,
//    CSRmreset       = 12'h782,
//    CSRmipi         = 12'h783,
//    CSRmiobase      = 12'h784
//} CSR deriving (Bits, Eq, FShow);
